module ins_mem(
input wire clk,
input wire rst,
input wire  [31:0] pc_in,
output wire [31:0] ins_out,
output wire [31:0] pc_out
);
wire [31:0] pc_increment;

endmodule;